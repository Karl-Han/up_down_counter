package test_pkg;
import env_pkg::*;

`include "test.sv"
endpackage