package env_pkg;
`include "transaction.sv"

`include "generator.sv"
`include "collector.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "environment.sv"
endpackage